library verilog;
use verilog.vl_types.all;
entity test_shepard is
end test_shepard;

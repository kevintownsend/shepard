library verilog;
use verilog.vl_types.all;
entity shepard is
    port(
        rst             : in     vl_logic;
        clk             : in     vl_logic;
        idle            : in     vl_logic;
        start           : in     vl_logic;
        stall           : out    vl_logic;
        aeId            : in     vl_logic_vector(1 downto 0);
        mc_req_ld_r0    : out    vl_logic;
        mc_req_vadr_r0  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_r0: in     vl_logic;
        mc_rsp_push_r0  : in     vl_logic;
        mc_rsp_stall_r0 : out    vl_logic;
        mc_rsp_data_r0  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_r1    : out    vl_logic;
        mc_req_vadr_r1  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_r1: in     vl_logic;
        mc_rsp_push_r1  : in     vl_logic;
        mc_rsp_stall_r1 : out    vl_logic;
        mc_rsp_data_r1  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_r2    : out    vl_logic;
        mc_req_vadr_r2  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_r2: in     vl_logic;
        mc_rsp_push_r2  : in     vl_logic;
        mc_rsp_stall_r2 : out    vl_logic;
        mc_rsp_data_r2  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_r3    : out    vl_logic;
        mc_req_vadr_r3  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_r3: in     vl_logic;
        mc_rsp_push_r3  : in     vl_logic;
        mc_rsp_stall_r3 : out    vl_logic;
        mc_rsp_data_r3  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_h0    : out    vl_logic;
        mc_req_vadr_h0  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_h0: in     vl_logic;
        mc_rsp_push_h0  : in     vl_logic;
        mc_rsp_stall_h0 : out    vl_logic;
        mc_rsp_data_h0  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_h1    : out    vl_logic;
        mc_req_vadr_h1  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_h1: in     vl_logic;
        mc_rsp_push_h1  : in     vl_logic;
        mc_rsp_stall_h1 : out    vl_logic;
        mc_rsp_data_h1  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_c0    : out    vl_logic;
        mc_req_vadr_c0  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_c0: in     vl_logic;
        mc_rsp_push_c0  : in     vl_logic;
        mc_rsp_stall_c0 : out    vl_logic;
        mc_rsp_data_c0  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_c1    : out    vl_logic;
        mc_req_vadr_c1  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_c1: in     vl_logic;
        mc_rsp_push_c1  : in     vl_logic;
        mc_rsp_stall_c1 : out    vl_logic;
        mc_rsp_data_c1  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_c2    : out    vl_logic;
        mc_req_vadr_c2  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_c2: in     vl_logic;
        mc_rsp_push_c2  : in     vl_logic;
        mc_rsp_stall_c2 : out    vl_logic;
        mc_rsp_data_c2  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_c3    : out    vl_logic;
        mc_req_vadr_c3  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_c3: in     vl_logic;
        mc_rsp_push_c3  : in     vl_logic;
        mc_rsp_stall_c3 : out    vl_logic;
        mc_rsp_data_c3  : in     vl_logic_vector(63 downto 0);
        mc_req_ld_c4    : out    vl_logic;
        mc_req_vadr_c4  : out    vl_logic_vector(47 downto 0);
        mc_rd_rq_stall_c4: in     vl_logic;
        mc_rsp_push_c4  : in     vl_logic;
        mc_rsp_stall_c4 : out    vl_logic;
        mc_rsp_data_c4  : in     vl_logic_vector(63 downto 0);
        mc_req_st_res   : out    vl_logic;
        mc_req_vadr_res : out    vl_logic_vector(47 downto 0);
        mc_req_data_res : out    vl_logic_vector(63 downto 0);
        mc_wr_rq_stall_res: in     vl_logic;
        hash_base       : in     vl_logic_vector(47 downto 0);
        hash_size       : in     vl_logic_vector(31 downto 0);
        ref_base        : in     vl_logic_vector(47 downto 0);
        read_base       : in     vl_logic_vector(47 downto 0);
        read_size       : in     vl_logic_vector(31 downto 0);
        res_base        : in     vl_logic_vector(47 downto 0)
    );
end shepard;

library verilog;
use verilog.vl_types.all;
entity hashTb is
end hashTb;
